module lcd(
	input rst,
	input clock,
	input [7:0] data
);

endmodule
