// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Wed Nov 04 16:27:59 2015

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    reset,clock,cond,
    output1);

    input reset;
    input clock;
    input cond;
    tri0 reset;
    tri0 cond;
    output output1;
    reg output1;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or cond)
    begin
        if (reset) begin
            reg_fstate <= state1;
            output1 <= 1'b0;
        end
        else begin
            output1 <= 1'b0;
            case (fstate)
                state1: begin
                    if ((cond == 1'b0))
                        reg_fstate <= state2;
                    else if ((cond == 1'b1))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    reg_fstate <= state3;
                end
                state3: begin
                    reg_fstate <= state4;

                    output1 <= 1'b1;
                end
                state4: begin
                    reg_fstate <= state5;
                end
                state5: begin
                    reg_fstate <= state1;

                    output1 <= 1'b0;
                end
                default: begin
                    output1 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
